module adder64 (cin,
    cout,
    a,
    b,
    s);
 input cin;
 output cout;
 input [63:0] a;
 input [63:0] b;
 output [63:0] s;

 wire c1;
 wire \Add1/c1 ;
 wire \Add1/c2 ;
 wire \Add1/c3 ;
 wire \Add1/Add1/c1 ;
 wire \Add1/Add1/Add1/_00_ ;
 wire \Add1/Add1/Add1/_01_ ;
 wire \Add1/Add1/Add1/_02_ ;
 wire \Add1/Add1/Add1/_03_ ;
 wire \Add1/Add1/Add1/_04_ ;
 wire \Add1/Add1/Add1/_05_ ;
 wire \Add1/Add1/Add1/_06_ ;
 wire \Add1/Add1/Add1/_07_ ;
 wire \Add1/Add1/Add1/_08_ ;
 wire \Add1/Add1/Add1/_09_ ;
 wire \Add1/Add1/Add1/_10_ ;
 wire \Add1/Add1/Add1/_11_ ;
 wire \Add1/Add1/Add1/_12_ ;
 wire \Add1/Add1/Add1/_13_ ;
 wire \Add1/Add1/Add1/_14_ ;
 wire \Add1/Add1/Add2/_00_ ;
 wire \Add1/Add1/Add2/_01_ ;
 wire \Add1/Add1/Add2/_02_ ;
 wire \Add1/Add1/Add2/_03_ ;
 wire \Add1/Add1/Add2/_04_ ;
 wire \Add1/Add1/Add2/_05_ ;
 wire \Add1/Add1/Add2/_06_ ;
 wire \Add1/Add1/Add2/_07_ ;
 wire \Add1/Add1/Add2/_08_ ;
 wire \Add1/Add1/Add2/_09_ ;
 wire \Add1/Add1/Add2/_10_ ;
 wire \Add1/Add1/Add2/_11_ ;
 wire \Add1/Add1/Add2/_12_ ;
 wire \Add1/Add1/Add2/_13_ ;
 wire \Add1/Add1/Add2/_14_ ;
 wire \Add1/Add2/c1 ;
 wire \Add1/Add2/Add1/_00_ ;
 wire \Add1/Add2/Add1/_01_ ;
 wire \Add1/Add2/Add1/_02_ ;
 wire \Add1/Add2/Add1/_03_ ;
 wire \Add1/Add2/Add1/_04_ ;
 wire \Add1/Add2/Add1/_05_ ;
 wire \Add1/Add2/Add1/_06_ ;
 wire \Add1/Add2/Add1/_07_ ;
 wire \Add1/Add2/Add1/_08_ ;
 wire \Add1/Add2/Add1/_09_ ;
 wire \Add1/Add2/Add1/_10_ ;
 wire \Add1/Add2/Add1/_11_ ;
 wire \Add1/Add2/Add1/_12_ ;
 wire \Add1/Add2/Add1/_13_ ;
 wire \Add1/Add2/Add1/_14_ ;
 wire \Add1/Add2/Add2/_00_ ;
 wire \Add1/Add2/Add2/_01_ ;
 wire \Add1/Add2/Add2/_02_ ;
 wire \Add1/Add2/Add2/_03_ ;
 wire \Add1/Add2/Add2/_04_ ;
 wire \Add1/Add2/Add2/_05_ ;
 wire \Add1/Add2/Add2/_06_ ;
 wire \Add1/Add2/Add2/_07_ ;
 wire \Add1/Add2/Add2/_08_ ;
 wire \Add1/Add2/Add2/_09_ ;
 wire \Add1/Add2/Add2/_10_ ;
 wire \Add1/Add2/Add2/_11_ ;
 wire \Add1/Add2/Add2/_12_ ;
 wire \Add1/Add2/Add2/_13_ ;
 wire \Add1/Add2/Add2/_14_ ;
 wire \Add1/Add3/c1 ;
 wire \Add1/Add3/Add1/_00_ ;
 wire \Add1/Add3/Add1/_01_ ;
 wire \Add1/Add3/Add1/_02_ ;
 wire \Add1/Add3/Add1/_03_ ;
 wire \Add1/Add3/Add1/_04_ ;
 wire \Add1/Add3/Add1/_05_ ;
 wire \Add1/Add3/Add1/_06_ ;
 wire \Add1/Add3/Add1/_07_ ;
 wire \Add1/Add3/Add1/_08_ ;
 wire \Add1/Add3/Add1/_09_ ;
 wire \Add1/Add3/Add1/_10_ ;
 wire \Add1/Add3/Add1/_11_ ;
 wire \Add1/Add3/Add1/_12_ ;
 wire \Add1/Add3/Add1/_13_ ;
 wire \Add1/Add3/Add1/_14_ ;
 wire \Add1/Add3/Add2/_00_ ;
 wire \Add1/Add3/Add2/_01_ ;
 wire \Add1/Add3/Add2/_02_ ;
 wire \Add1/Add3/Add2/_03_ ;
 wire \Add1/Add3/Add2/_04_ ;
 wire \Add1/Add3/Add2/_05_ ;
 wire \Add1/Add3/Add2/_06_ ;
 wire \Add1/Add3/Add2/_07_ ;
 wire \Add1/Add3/Add2/_08_ ;
 wire \Add1/Add3/Add2/_09_ ;
 wire \Add1/Add3/Add2/_10_ ;
 wire \Add1/Add3/Add2/_11_ ;
 wire \Add1/Add3/Add2/_12_ ;
 wire \Add1/Add3/Add2/_13_ ;
 wire \Add1/Add3/Add2/_14_ ;
 wire \Add1/Add4/c1 ;
 wire \Add1/Add4/Add1/_00_ ;
 wire \Add1/Add4/Add1/_01_ ;
 wire \Add1/Add4/Add1/_02_ ;
 wire \Add1/Add4/Add1/_03_ ;
 wire \Add1/Add4/Add1/_04_ ;
 wire \Add1/Add4/Add1/_05_ ;
 wire \Add1/Add4/Add1/_06_ ;
 wire \Add1/Add4/Add1/_07_ ;
 wire \Add1/Add4/Add1/_08_ ;
 wire \Add1/Add4/Add1/_09_ ;
 wire \Add1/Add4/Add1/_10_ ;
 wire \Add1/Add4/Add1/_11_ ;
 wire \Add1/Add4/Add1/_12_ ;
 wire \Add1/Add4/Add1/_13_ ;
 wire \Add1/Add4/Add1/_14_ ;
 wire \Add1/Add4/Add2/_00_ ;
 wire \Add1/Add4/Add2/_01_ ;
 wire \Add1/Add4/Add2/_02_ ;
 wire \Add1/Add4/Add2/_03_ ;
 wire \Add1/Add4/Add2/_04_ ;
 wire \Add1/Add4/Add2/_05_ ;
 wire \Add1/Add4/Add2/_06_ ;
 wire \Add1/Add4/Add2/_07_ ;
 wire \Add1/Add4/Add2/_08_ ;
 wire \Add1/Add4/Add2/_09_ ;
 wire \Add1/Add4/Add2/_10_ ;
 wire \Add1/Add4/Add2/_11_ ;
 wire \Add1/Add4/Add2/_12_ ;
 wire \Add1/Add4/Add2/_13_ ;
 wire \Add1/Add4/Add2/_14_ ;
 wire \Add2/c1 ;
 wire \Add2/c2 ;
 wire \Add2/c3 ;
 wire \Add2/Add1/c1 ;
 wire \Add2/Add1/Add1/_00_ ;
 wire \Add2/Add1/Add1/_01_ ;
 wire \Add2/Add1/Add1/_02_ ;
 wire \Add2/Add1/Add1/_03_ ;
 wire \Add2/Add1/Add1/_04_ ;
 wire \Add2/Add1/Add1/_05_ ;
 wire \Add2/Add1/Add1/_06_ ;
 wire \Add2/Add1/Add1/_07_ ;
 wire \Add2/Add1/Add1/_08_ ;
 wire \Add2/Add1/Add1/_09_ ;
 wire \Add2/Add1/Add1/_10_ ;
 wire \Add2/Add1/Add1/_11_ ;
 wire \Add2/Add1/Add1/_12_ ;
 wire \Add2/Add1/Add1/_13_ ;
 wire \Add2/Add1/Add1/_14_ ;
 wire \Add2/Add1/Add2/_00_ ;
 wire \Add2/Add1/Add2/_01_ ;
 wire \Add2/Add1/Add2/_02_ ;
 wire \Add2/Add1/Add2/_03_ ;
 wire \Add2/Add1/Add2/_04_ ;
 wire \Add2/Add1/Add2/_05_ ;
 wire \Add2/Add1/Add2/_06_ ;
 wire \Add2/Add1/Add2/_07_ ;
 wire \Add2/Add1/Add2/_08_ ;
 wire \Add2/Add1/Add2/_09_ ;
 wire \Add2/Add1/Add2/_10_ ;
 wire \Add2/Add1/Add2/_11_ ;
 wire \Add2/Add1/Add2/_12_ ;
 wire \Add2/Add1/Add2/_13_ ;
 wire \Add2/Add1/Add2/_14_ ;
 wire \Add2/Add2/c1 ;
 wire \Add2/Add2/Add1/_00_ ;
 wire \Add2/Add2/Add1/_01_ ;
 wire \Add2/Add2/Add1/_02_ ;
 wire \Add2/Add2/Add1/_03_ ;
 wire \Add2/Add2/Add1/_04_ ;
 wire \Add2/Add2/Add1/_05_ ;
 wire \Add2/Add2/Add1/_06_ ;
 wire \Add2/Add2/Add1/_07_ ;
 wire \Add2/Add2/Add1/_08_ ;
 wire \Add2/Add2/Add1/_09_ ;
 wire \Add2/Add2/Add1/_10_ ;
 wire \Add2/Add2/Add1/_11_ ;
 wire \Add2/Add2/Add1/_12_ ;
 wire \Add2/Add2/Add1/_13_ ;
 wire \Add2/Add2/Add1/_14_ ;
 wire \Add2/Add2/Add2/_00_ ;
 wire \Add2/Add2/Add2/_01_ ;
 wire \Add2/Add2/Add2/_02_ ;
 wire \Add2/Add2/Add2/_03_ ;
 wire \Add2/Add2/Add2/_04_ ;
 wire \Add2/Add2/Add2/_05_ ;
 wire \Add2/Add2/Add2/_06_ ;
 wire \Add2/Add2/Add2/_07_ ;
 wire \Add2/Add2/Add2/_08_ ;
 wire \Add2/Add2/Add2/_09_ ;
 wire \Add2/Add2/Add2/_10_ ;
 wire \Add2/Add2/Add2/_11_ ;
 wire \Add2/Add2/Add2/_12_ ;
 wire \Add2/Add2/Add2/_13_ ;
 wire \Add2/Add2/Add2/_14_ ;
 wire \Add2/Add3/c1 ;
 wire \Add2/Add3/Add1/_00_ ;
 wire \Add2/Add3/Add1/_01_ ;
 wire \Add2/Add3/Add1/_02_ ;
 wire \Add2/Add3/Add1/_03_ ;
 wire \Add2/Add3/Add1/_04_ ;
 wire \Add2/Add3/Add1/_05_ ;
 wire \Add2/Add3/Add1/_06_ ;
 wire \Add2/Add3/Add1/_07_ ;
 wire \Add2/Add3/Add1/_08_ ;
 wire \Add2/Add3/Add1/_09_ ;
 wire \Add2/Add3/Add1/_10_ ;
 wire \Add2/Add3/Add1/_11_ ;
 wire \Add2/Add3/Add1/_12_ ;
 wire \Add2/Add3/Add1/_13_ ;
 wire \Add2/Add3/Add1/_14_ ;
 wire \Add2/Add3/Add2/_00_ ;
 wire \Add2/Add3/Add2/_01_ ;
 wire \Add2/Add3/Add2/_02_ ;
 wire \Add2/Add3/Add2/_03_ ;
 wire \Add2/Add3/Add2/_04_ ;
 wire \Add2/Add3/Add2/_05_ ;
 wire \Add2/Add3/Add2/_06_ ;
 wire \Add2/Add3/Add2/_07_ ;
 wire \Add2/Add3/Add2/_08_ ;
 wire \Add2/Add3/Add2/_09_ ;
 wire \Add2/Add3/Add2/_10_ ;
 wire \Add2/Add3/Add2/_11_ ;
 wire \Add2/Add3/Add2/_12_ ;
 wire \Add2/Add3/Add2/_13_ ;
 wire \Add2/Add3/Add2/_14_ ;
 wire \Add2/Add4/c1 ;
 wire \Add2/Add4/Add1/_00_ ;
 wire \Add2/Add4/Add1/_01_ ;
 wire \Add2/Add4/Add1/_02_ ;
 wire \Add2/Add4/Add1/_03_ ;
 wire \Add2/Add4/Add1/_04_ ;
 wire \Add2/Add4/Add1/_05_ ;
 wire \Add2/Add4/Add1/_06_ ;
 wire \Add2/Add4/Add1/_07_ ;
 wire \Add2/Add4/Add1/_08_ ;
 wire \Add2/Add4/Add1/_09_ ;
 wire \Add2/Add4/Add1/_10_ ;
 wire \Add2/Add4/Add1/_11_ ;
 wire \Add2/Add4/Add1/_12_ ;
 wire \Add2/Add4/Add1/_13_ ;
 wire \Add2/Add4/Add1/_14_ ;
 wire \Add2/Add4/Add2/_00_ ;
 wire \Add2/Add4/Add2/_01_ ;
 wire \Add2/Add4/Add2/_02_ ;
 wire \Add2/Add4/Add2/_03_ ;
 wire \Add2/Add4/Add2/_04_ ;
 wire \Add2/Add4/Add2/_05_ ;
 wire \Add2/Add4/Add2/_06_ ;
 wire \Add2/Add4/Add2/_07_ ;
 wire \Add2/Add4/Add2/_08_ ;
 wire \Add2/Add4/Add2/_09_ ;
 wire \Add2/Add4/Add2/_10_ ;
 wire \Add2/Add4/Add2/_11_ ;
 wire \Add2/Add4/Add2/_12_ ;
 wire \Add2/Add4/Add2/_13_ ;
 wire \Add2/Add4/Add2/_14_ ;

 NAND2_X1 \Add1/Add1/Add1/_15_  (.A1(a[3]),
    .A2(b[3]),
    .ZN(\Add1/Add1/Add1/_00_ ));
 AND2_X1 \Add1/Add1/Add1/_16_  (.A1(a[2]),
    .A2(b[2]),
    .ZN(\Add1/Add1/Add1/_01_ ));
 NAND2_X1 \Add1/Add1/Add1/_17_  (.A1(a[1]),
    .A2(b[1]),
    .ZN(\Add1/Add1/Add1/_02_ ));
 AND2_X1 \Add1/Add1/Add1/_18_  (.A1(a[0]),
    .A2(b[0]),
    .ZN(\Add1/Add1/Add1/_03_ ));
 OR2_X1 \Add1/Add1/Add1/_19_  (.A1(a[0]),
    .A2(b[0]),
    .ZN(\Add1/Add1/Add1/_04_ ));
 XNOR2_X1 \Add1/Add1/Add1/_20_  (.A(a[0]),
    .B(b[0]),
    .ZN(\Add1/Add1/Add1/_05_ ));
 AOI21_X2 \Add1/Add1/Add1/_21_  (.A(\Add1/Add1/Add1/_03_ ),
    .B1(\Add1/Add1/Add1/_04_ ),
    .B2(cin),
    .ZN(\Add1/Add1/Add1/_06_ ));
 NOR2_X1 \Add1/Add1/Add1/_22_  (.A1(a[1]),
    .A2(b[1]),
    .ZN(\Add1/Add1/Add1/_07_ ));
 XOR2_X1 \Add1/Add1/Add1/_23_  (.A(a[1]),
    .B(b[1]),
    .Z(\Add1/Add1/Add1/_08_ ));
 OAI21_X2 \Add1/Add1/Add1/_24_  (.A(\Add1/Add1/Add1/_02_ ),
    .B1(\Add1/Add1/Add1/_06_ ),
    .B2(\Add1/Add1/Add1/_07_ ),
    .ZN(\Add1/Add1/Add1/_09_ ));
 OR2_X1 \Add1/Add1/Add1/_25_  (.A1(a[2]),
    .A2(b[2]),
    .ZN(\Add1/Add1/Add1/_10_ ));
 XNOR2_X1 \Add1/Add1/Add1/_26_  (.A(a[2]),
    .B(b[2]),
    .ZN(\Add1/Add1/Add1/_11_ ));
 AOI21_X2 \Add1/Add1/Add1/_27_  (.A(\Add1/Add1/Add1/_01_ ),
    .B1(\Add1/Add1/Add1/_09_ ),
    .B2(\Add1/Add1/Add1/_10_ ),
    .ZN(\Add1/Add1/Add1/_12_ ));
 NOR2_X1 \Add1/Add1/Add1/_28_  (.A1(a[3]),
    .A2(b[3]),
    .ZN(\Add1/Add1/Add1/_13_ ));
 XOR2_X1 \Add1/Add1/Add1/_29_  (.A(a[3]),
    .B(b[3]),
    .Z(\Add1/Add1/Add1/_14_ ));
 OAI21_X2 \Add1/Add1/Add1/_30_  (.A(\Add1/Add1/Add1/_00_ ),
    .B1(\Add1/Add1/Add1/_12_ ),
    .B2(\Add1/Add1/Add1/_13_ ),
    .ZN(\Add1/Add1/c1 ));
 XNOR2_X1 \Add1/Add1/Add1/_31_  (.A(cin),
    .B(\Add1/Add1/Add1/_05_ ),
    .ZN(s[0]));
 XNOR2_X1 \Add1/Add1/Add1/_32_  (.A(\Add1/Add1/Add1/_06_ ),
    .B(\Add1/Add1/Add1/_08_ ),
    .ZN(s[1]));
 XNOR2_X1 \Add1/Add1/Add1/_33_  (.A(\Add1/Add1/Add1/_09_ ),
    .B(\Add1/Add1/Add1/_11_ ),
    .ZN(s[2]));
 XNOR2_X1 \Add1/Add1/Add1/_34_  (.A(\Add1/Add1/Add1/_12_ ),
    .B(\Add1/Add1/Add1/_14_ ),
    .ZN(s[3]));
 NAND2_X1 \Add1/Add1/Add2/_15_  (.A1(a[7]),
    .A2(b[7]),
    .ZN(\Add1/Add1/Add2/_00_ ));
 AND2_X1 \Add1/Add1/Add2/_16_  (.A1(a[6]),
    .A2(b[6]),
    .ZN(\Add1/Add1/Add2/_01_ ));
 NAND2_X1 \Add1/Add1/Add2/_17_  (.A1(a[5]),
    .A2(b[5]),
    .ZN(\Add1/Add1/Add2/_02_ ));
 AND2_X1 \Add1/Add1/Add2/_18_  (.A1(a[4]),
    .A2(b[4]),
    .ZN(\Add1/Add1/Add2/_03_ ));
 OR2_X1 \Add1/Add1/Add2/_19_  (.A1(a[4]),
    .A2(b[4]),
    .ZN(\Add1/Add1/Add2/_04_ ));
 XNOR2_X1 \Add1/Add1/Add2/_20_  (.A(a[4]),
    .B(b[4]),
    .ZN(\Add1/Add1/Add2/_05_ ));
 AOI21_X4 \Add1/Add1/Add2/_21_  (.A(\Add1/Add1/Add2/_03_ ),
    .B1(\Add1/Add1/Add2/_04_ ),
    .B2(\Add1/Add1/c1 ),
    .ZN(\Add1/Add1/Add2/_06_ ));
 NOR2_X1 \Add1/Add1/Add2/_22_  (.A1(a[5]),
    .A2(b[5]),
    .ZN(\Add1/Add1/Add2/_07_ ));
 XOR2_X1 \Add1/Add1/Add2/_23_  (.A(a[5]),
    .B(b[5]),
    .Z(\Add1/Add1/Add2/_08_ ));
 OAI21_X2 \Add1/Add1/Add2/_24_  (.A(\Add1/Add1/Add2/_02_ ),
    .B1(\Add1/Add1/Add2/_06_ ),
    .B2(\Add1/Add1/Add2/_07_ ),
    .ZN(\Add1/Add1/Add2/_09_ ));
 OR2_X1 \Add1/Add1/Add2/_25_  (.A1(a[6]),
    .A2(b[6]),
    .ZN(\Add1/Add1/Add2/_10_ ));
 XNOR2_X1 \Add1/Add1/Add2/_26_  (.A(a[6]),
    .B(b[6]),
    .ZN(\Add1/Add1/Add2/_11_ ));
 AOI21_X4 \Add1/Add1/Add2/_27_  (.A(\Add1/Add1/Add2/_01_ ),
    .B1(\Add1/Add1/Add2/_09_ ),
    .B2(\Add1/Add1/Add2/_10_ ),
    .ZN(\Add1/Add1/Add2/_12_ ));
 NOR2_X1 \Add1/Add1/Add2/_28_  (.A1(a[7]),
    .A2(b[7]),
    .ZN(\Add1/Add1/Add2/_13_ ));
 XOR2_X1 \Add1/Add1/Add2/_29_  (.A(a[7]),
    .B(b[7]),
    .Z(\Add1/Add1/Add2/_14_ ));
 OAI21_X1 \Add1/Add1/Add2/_30_  (.A(\Add1/Add1/Add2/_00_ ),
    .B1(\Add1/Add1/Add2/_12_ ),
    .B2(\Add1/Add1/Add2/_13_ ),
    .ZN(\Add1/c1 ));
 XNOR2_X1 \Add1/Add1/Add2/_31_  (.A(\Add1/Add1/c1 ),
    .B(\Add1/Add1/Add2/_05_ ),
    .ZN(s[4]));
 XNOR2_X1 \Add1/Add1/Add2/_32_  (.A(\Add1/Add1/Add2/_06_ ),
    .B(\Add1/Add1/Add2/_08_ ),
    .ZN(s[5]));
 XNOR2_X1 \Add1/Add1/Add2/_33_  (.A(\Add1/Add1/Add2/_09_ ),
    .B(\Add1/Add1/Add2/_11_ ),
    .ZN(s[6]));
 XNOR2_X1 \Add1/Add1/Add2/_34_  (.A(\Add1/Add1/Add2/_12_ ),
    .B(\Add1/Add1/Add2/_14_ ),
    .ZN(s[7]));
 NAND2_X1 \Add1/Add2/Add1/_15_  (.A1(a[11]),
    .A2(b[11]),
    .ZN(\Add1/Add2/Add1/_00_ ));
 AND2_X1 \Add1/Add2/Add1/_16_  (.A1(a[10]),
    .A2(b[10]),
    .ZN(\Add1/Add2/Add1/_01_ ));
 NAND2_X1 \Add1/Add2/Add1/_17_  (.A1(a[9]),
    .A2(b[9]),
    .ZN(\Add1/Add2/Add1/_02_ ));
 AND2_X1 \Add1/Add2/Add1/_18_  (.A1(a[8]),
    .A2(b[8]),
    .ZN(\Add1/Add2/Add1/_03_ ));
 OR2_X1 \Add1/Add2/Add1/_19_  (.A1(a[8]),
    .A2(b[8]),
    .ZN(\Add1/Add2/Add1/_04_ ));
 XNOR2_X1 \Add1/Add2/Add1/_20_  (.A(a[8]),
    .B(b[8]),
    .ZN(\Add1/Add2/Add1/_05_ ));
 AOI21_X1 \Add1/Add2/Add1/_21_  (.A(\Add1/Add2/Add1/_03_ ),
    .B1(\Add1/Add2/Add1/_04_ ),
    .B2(\Add1/c1 ),
    .ZN(\Add1/Add2/Add1/_06_ ));
 NOR2_X1 \Add1/Add2/Add1/_22_  (.A1(a[9]),
    .A2(b[9]),
    .ZN(\Add1/Add2/Add1/_07_ ));
 XOR2_X1 \Add1/Add2/Add1/_23_  (.A(a[9]),
    .B(b[9]),
    .Z(\Add1/Add2/Add1/_08_ ));
 OAI21_X1 \Add1/Add2/Add1/_24_  (.A(\Add1/Add2/Add1/_02_ ),
    .B1(\Add1/Add2/Add1/_06_ ),
    .B2(\Add1/Add2/Add1/_07_ ),
    .ZN(\Add1/Add2/Add1/_09_ ));
 OR2_X1 \Add1/Add2/Add1/_25_  (.A1(a[10]),
    .A2(b[10]),
    .ZN(\Add1/Add2/Add1/_10_ ));
 XNOR2_X1 \Add1/Add2/Add1/_26_  (.A(a[10]),
    .B(b[10]),
    .ZN(\Add1/Add2/Add1/_11_ ));
 AOI21_X1 \Add1/Add2/Add1/_27_  (.A(\Add1/Add2/Add1/_01_ ),
    .B1(\Add1/Add2/Add1/_09_ ),
    .B2(\Add1/Add2/Add1/_10_ ),
    .ZN(\Add1/Add2/Add1/_12_ ));
 NOR2_X1 \Add1/Add2/Add1/_28_  (.A1(a[11]),
    .A2(b[11]),
    .ZN(\Add1/Add2/Add1/_13_ ));
 XOR2_X1 \Add1/Add2/Add1/_29_  (.A(a[11]),
    .B(b[11]),
    .Z(\Add1/Add2/Add1/_14_ ));
 OAI21_X1 \Add1/Add2/Add1/_30_  (.A(\Add1/Add2/Add1/_00_ ),
    .B1(\Add1/Add2/Add1/_12_ ),
    .B2(\Add1/Add2/Add1/_13_ ),
    .ZN(\Add1/Add2/c1 ));
 XNOR2_X1 \Add1/Add2/Add1/_31_  (.A(\Add1/c1 ),
    .B(\Add1/Add2/Add1/_05_ ),
    .ZN(s[8]));
 XNOR2_X1 \Add1/Add2/Add1/_32_  (.A(\Add1/Add2/Add1/_06_ ),
    .B(\Add1/Add2/Add1/_08_ ),
    .ZN(s[9]));
 XNOR2_X1 \Add1/Add2/Add1/_33_  (.A(\Add1/Add2/Add1/_09_ ),
    .B(\Add1/Add2/Add1/_11_ ),
    .ZN(s[10]));
 XNOR2_X1 \Add1/Add2/Add1/_34_  (.A(\Add1/Add2/Add1/_12_ ),
    .B(\Add1/Add2/Add1/_14_ ),
    .ZN(s[11]));
 NAND2_X1 \Add1/Add2/Add2/_15_  (.A1(a[15]),
    .A2(b[15]),
    .ZN(\Add1/Add2/Add2/_00_ ));
 AND2_X1 \Add1/Add2/Add2/_16_  (.A1(a[14]),
    .A2(b[14]),
    .ZN(\Add1/Add2/Add2/_01_ ));
 NAND2_X1 \Add1/Add2/Add2/_17_  (.A1(a[13]),
    .A2(b[13]),
    .ZN(\Add1/Add2/Add2/_02_ ));
 AND2_X1 \Add1/Add2/Add2/_18_  (.A1(a[12]),
    .A2(b[12]),
    .ZN(\Add1/Add2/Add2/_03_ ));
 OR2_X1 \Add1/Add2/Add2/_19_  (.A1(a[12]),
    .A2(b[12]),
    .ZN(\Add1/Add2/Add2/_04_ ));
 XNOR2_X1 \Add1/Add2/Add2/_20_  (.A(a[12]),
    .B(b[12]),
    .ZN(\Add1/Add2/Add2/_05_ ));
 AOI21_X2 \Add1/Add2/Add2/_21_  (.A(\Add1/Add2/Add2/_03_ ),
    .B1(\Add1/Add2/Add2/_04_ ),
    .B2(\Add1/Add2/c1 ),
    .ZN(\Add1/Add2/Add2/_06_ ));
 NOR2_X1 \Add1/Add2/Add2/_22_  (.A1(a[13]),
    .A2(b[13]),
    .ZN(\Add1/Add2/Add2/_07_ ));
 XOR2_X1 \Add1/Add2/Add2/_23_  (.A(a[13]),
    .B(b[13]),
    .Z(\Add1/Add2/Add2/_08_ ));
 OAI21_X2 \Add1/Add2/Add2/_24_  (.A(\Add1/Add2/Add2/_02_ ),
    .B1(\Add1/Add2/Add2/_06_ ),
    .B2(\Add1/Add2/Add2/_07_ ),
    .ZN(\Add1/Add2/Add2/_09_ ));
 OR2_X1 \Add1/Add2/Add2/_25_  (.A1(a[14]),
    .A2(b[14]),
    .ZN(\Add1/Add2/Add2/_10_ ));
 XNOR2_X1 \Add1/Add2/Add2/_26_  (.A(a[14]),
    .B(b[14]),
    .ZN(\Add1/Add2/Add2/_11_ ));
 AOI21_X2 \Add1/Add2/Add2/_27_  (.A(\Add1/Add2/Add2/_01_ ),
    .B1(\Add1/Add2/Add2/_09_ ),
    .B2(\Add1/Add2/Add2/_10_ ),
    .ZN(\Add1/Add2/Add2/_12_ ));
 NOR2_X1 \Add1/Add2/Add2/_28_  (.A1(a[15]),
    .A2(b[15]),
    .ZN(\Add1/Add2/Add2/_13_ ));
 XOR2_X1 \Add1/Add2/Add2/_29_  (.A(a[15]),
    .B(b[15]),
    .Z(\Add1/Add2/Add2/_14_ ));
 OAI21_X4 \Add1/Add2/Add2/_30_  (.A(\Add1/Add2/Add2/_00_ ),
    .B1(\Add1/Add2/Add2/_12_ ),
    .B2(\Add1/Add2/Add2/_13_ ),
    .ZN(\Add1/c2 ));
 XNOR2_X1 \Add1/Add2/Add2/_31_  (.A(\Add1/Add2/c1 ),
    .B(\Add1/Add2/Add2/_05_ ),
    .ZN(s[12]));
 XNOR2_X1 \Add1/Add2/Add2/_32_  (.A(\Add1/Add2/Add2/_06_ ),
    .B(\Add1/Add2/Add2/_08_ ),
    .ZN(s[13]));
 XNOR2_X1 \Add1/Add2/Add2/_33_  (.A(\Add1/Add2/Add2/_09_ ),
    .B(\Add1/Add2/Add2/_11_ ),
    .ZN(s[14]));
 XNOR2_X1 \Add1/Add2/Add2/_34_  (.A(\Add1/Add2/Add2/_12_ ),
    .B(\Add1/Add2/Add2/_14_ ),
    .ZN(s[15]));
 NAND2_X1 \Add1/Add3/Add1/_15_  (.A1(a[19]),
    .A2(b[19]),
    .ZN(\Add1/Add3/Add1/_00_ ));
 AND2_X1 \Add1/Add3/Add1/_16_  (.A1(a[18]),
    .A2(b[18]),
    .ZN(\Add1/Add3/Add1/_01_ ));
 NAND2_X1 \Add1/Add3/Add1/_17_  (.A1(a[17]),
    .A2(b[17]),
    .ZN(\Add1/Add3/Add1/_02_ ));
 AND2_X1 \Add1/Add3/Add1/_18_  (.A1(a[16]),
    .A2(b[16]),
    .ZN(\Add1/Add3/Add1/_03_ ));
 OR2_X1 \Add1/Add3/Add1/_19_  (.A1(a[16]),
    .A2(b[16]),
    .ZN(\Add1/Add3/Add1/_04_ ));
 XNOR2_X1 \Add1/Add3/Add1/_20_  (.A(a[16]),
    .B(b[16]),
    .ZN(\Add1/Add3/Add1/_05_ ));
 AOI21_X2 \Add1/Add3/Add1/_21_  (.A(\Add1/Add3/Add1/_03_ ),
    .B1(\Add1/Add3/Add1/_04_ ),
    .B2(\Add1/c2 ),
    .ZN(\Add1/Add3/Add1/_06_ ));
 NOR2_X1 \Add1/Add3/Add1/_22_  (.A1(a[17]),
    .A2(b[17]),
    .ZN(\Add1/Add3/Add1/_07_ ));
 XOR2_X1 \Add1/Add3/Add1/_23_  (.A(a[17]),
    .B(b[17]),
    .Z(\Add1/Add3/Add1/_08_ ));
 OAI21_X2 \Add1/Add3/Add1/_24_  (.A(\Add1/Add3/Add1/_02_ ),
    .B1(\Add1/Add3/Add1/_06_ ),
    .B2(\Add1/Add3/Add1/_07_ ),
    .ZN(\Add1/Add3/Add1/_09_ ));
 OR2_X1 \Add1/Add3/Add1/_25_  (.A1(a[18]),
    .A2(b[18]),
    .ZN(\Add1/Add3/Add1/_10_ ));
 XNOR2_X1 \Add1/Add3/Add1/_26_  (.A(a[18]),
    .B(b[18]),
    .ZN(\Add1/Add3/Add1/_11_ ));
 AOI21_X2 \Add1/Add3/Add1/_27_  (.A(\Add1/Add3/Add1/_01_ ),
    .B1(\Add1/Add3/Add1/_09_ ),
    .B2(\Add1/Add3/Add1/_10_ ),
    .ZN(\Add1/Add3/Add1/_12_ ));
 NOR2_X1 \Add1/Add3/Add1/_28_  (.A1(a[19]),
    .A2(b[19]),
    .ZN(\Add1/Add3/Add1/_13_ ));
 XOR2_X1 \Add1/Add3/Add1/_29_  (.A(a[19]),
    .B(b[19]),
    .Z(\Add1/Add3/Add1/_14_ ));
 OAI21_X4 \Add1/Add3/Add1/_30_  (.A(\Add1/Add3/Add1/_00_ ),
    .B1(\Add1/Add3/Add1/_12_ ),
    .B2(\Add1/Add3/Add1/_13_ ),
    .ZN(\Add1/Add3/c1 ));
 XNOR2_X1 \Add1/Add3/Add1/_31_  (.A(\Add1/c2 ),
    .B(\Add1/Add3/Add1/_05_ ),
    .ZN(s[16]));
 XNOR2_X1 \Add1/Add3/Add1/_32_  (.A(\Add1/Add3/Add1/_06_ ),
    .B(\Add1/Add3/Add1/_08_ ),
    .ZN(s[17]));
 XNOR2_X1 \Add1/Add3/Add1/_33_  (.A(\Add1/Add3/Add1/_09_ ),
    .B(\Add1/Add3/Add1/_11_ ),
    .ZN(s[18]));
 XNOR2_X1 \Add1/Add3/Add1/_34_  (.A(\Add1/Add3/Add1/_12_ ),
    .B(\Add1/Add3/Add1/_14_ ),
    .ZN(s[19]));
 NAND2_X1 \Add1/Add3/Add2/_15_  (.A1(a[23]),
    .A2(b[23]),
    .ZN(\Add1/Add3/Add2/_00_ ));
 AND2_X1 \Add1/Add3/Add2/_16_  (.A1(a[22]),
    .A2(b[22]),
    .ZN(\Add1/Add3/Add2/_01_ ));
 NAND2_X1 \Add1/Add3/Add2/_17_  (.A1(a[21]),
    .A2(b[21]),
    .ZN(\Add1/Add3/Add2/_02_ ));
 AND2_X1 \Add1/Add3/Add2/_18_  (.A1(a[20]),
    .A2(b[20]),
    .ZN(\Add1/Add3/Add2/_03_ ));
 OR2_X1 \Add1/Add3/Add2/_19_  (.A1(a[20]),
    .A2(b[20]),
    .ZN(\Add1/Add3/Add2/_04_ ));
 XNOR2_X1 \Add1/Add3/Add2/_20_  (.A(a[20]),
    .B(b[20]),
    .ZN(\Add1/Add3/Add2/_05_ ));
 AOI21_X4 \Add1/Add3/Add2/_21_  (.A(\Add1/Add3/Add2/_03_ ),
    .B1(\Add1/Add3/Add2/_04_ ),
    .B2(\Add1/Add3/c1 ),
    .ZN(\Add1/Add3/Add2/_06_ ));
 NOR2_X1 \Add1/Add3/Add2/_22_  (.A1(a[21]),
    .A2(b[21]),
    .ZN(\Add1/Add3/Add2/_07_ ));
 XOR2_X1 \Add1/Add3/Add2/_23_  (.A(a[21]),
    .B(b[21]),
    .Z(\Add1/Add3/Add2/_08_ ));
 OAI21_X1 \Add1/Add3/Add2/_24_  (.A(\Add1/Add3/Add2/_02_ ),
    .B1(\Add1/Add3/Add2/_06_ ),
    .B2(\Add1/Add3/Add2/_07_ ),
    .ZN(\Add1/Add3/Add2/_09_ ));
 OR2_X1 \Add1/Add3/Add2/_25_  (.A1(a[22]),
    .A2(b[22]),
    .ZN(\Add1/Add3/Add2/_10_ ));
 XNOR2_X1 \Add1/Add3/Add2/_26_  (.A(a[22]),
    .B(b[22]),
    .ZN(\Add1/Add3/Add2/_11_ ));
 AOI21_X2 \Add1/Add3/Add2/_27_  (.A(\Add1/Add3/Add2/_01_ ),
    .B1(\Add1/Add3/Add2/_09_ ),
    .B2(\Add1/Add3/Add2/_10_ ),
    .ZN(\Add1/Add3/Add2/_12_ ));
 NOR2_X1 \Add1/Add3/Add2/_28_  (.A1(a[23]),
    .A2(b[23]),
    .ZN(\Add1/Add3/Add2/_13_ ));
 XOR2_X1 \Add1/Add3/Add2/_29_  (.A(a[23]),
    .B(b[23]),
    .Z(\Add1/Add3/Add2/_14_ ));
 OAI21_X2 \Add1/Add3/Add2/_30_  (.A(\Add1/Add3/Add2/_00_ ),
    .B1(\Add1/Add3/Add2/_12_ ),
    .B2(\Add1/Add3/Add2/_13_ ),
    .ZN(\Add1/c3 ));
 XNOR2_X1 \Add1/Add3/Add2/_31_  (.A(\Add1/Add3/c1 ),
    .B(\Add1/Add3/Add2/_05_ ),
    .ZN(s[20]));
 XNOR2_X1 \Add1/Add3/Add2/_32_  (.A(\Add1/Add3/Add2/_06_ ),
    .B(\Add1/Add3/Add2/_08_ ),
    .ZN(s[21]));
 XNOR2_X1 \Add1/Add3/Add2/_33_  (.A(\Add1/Add3/Add2/_09_ ),
    .B(\Add1/Add3/Add2/_11_ ),
    .ZN(s[22]));
 XNOR2_X1 \Add1/Add3/Add2/_34_  (.A(\Add1/Add3/Add2/_12_ ),
    .B(\Add1/Add3/Add2/_14_ ),
    .ZN(s[23]));
 NAND2_X1 \Add1/Add4/Add1/_15_  (.A1(a[27]),
    .A2(b[27]),
    .ZN(\Add1/Add4/Add1/_00_ ));
 AND2_X1 \Add1/Add4/Add1/_16_  (.A1(a[26]),
    .A2(b[26]),
    .ZN(\Add1/Add4/Add1/_01_ ));
 NAND2_X1 \Add1/Add4/Add1/_17_  (.A1(a[25]),
    .A2(b[25]),
    .ZN(\Add1/Add4/Add1/_02_ ));
 AND2_X1 \Add1/Add4/Add1/_18_  (.A1(a[24]),
    .A2(b[24]),
    .ZN(\Add1/Add4/Add1/_03_ ));
 OR2_X1 \Add1/Add4/Add1/_19_  (.A1(a[24]),
    .A2(b[24]),
    .ZN(\Add1/Add4/Add1/_04_ ));
 XNOR2_X1 \Add1/Add4/Add1/_20_  (.A(a[24]),
    .B(b[24]),
    .ZN(\Add1/Add4/Add1/_05_ ));
 AOI21_X4 \Add1/Add4/Add1/_21_  (.A(\Add1/Add4/Add1/_03_ ),
    .B1(\Add1/Add4/Add1/_04_ ),
    .B2(\Add1/c3 ),
    .ZN(\Add1/Add4/Add1/_06_ ));
 NOR2_X1 \Add1/Add4/Add1/_22_  (.A1(a[25]),
    .A2(b[25]),
    .ZN(\Add1/Add4/Add1/_07_ ));
 XOR2_X1 \Add1/Add4/Add1/_23_  (.A(a[25]),
    .B(b[25]),
    .Z(\Add1/Add4/Add1/_08_ ));
 OAI21_X2 \Add1/Add4/Add1/_24_  (.A(\Add1/Add4/Add1/_02_ ),
    .B1(\Add1/Add4/Add1/_06_ ),
    .B2(\Add1/Add4/Add1/_07_ ),
    .ZN(\Add1/Add4/Add1/_09_ ));
 OR2_X1 \Add1/Add4/Add1/_25_  (.A1(a[26]),
    .A2(b[26]),
    .ZN(\Add1/Add4/Add1/_10_ ));
 XNOR2_X1 \Add1/Add4/Add1/_26_  (.A(a[26]),
    .B(b[26]),
    .ZN(\Add1/Add4/Add1/_11_ ));
 AOI21_X4 \Add1/Add4/Add1/_27_  (.A(\Add1/Add4/Add1/_01_ ),
    .B1(\Add1/Add4/Add1/_09_ ),
    .B2(\Add1/Add4/Add1/_10_ ),
    .ZN(\Add1/Add4/Add1/_12_ ));
 NOR2_X1 \Add1/Add4/Add1/_28_  (.A1(a[27]),
    .A2(b[27]),
    .ZN(\Add1/Add4/Add1/_13_ ));
 XOR2_X1 \Add1/Add4/Add1/_29_  (.A(a[27]),
    .B(b[27]),
    .Z(\Add1/Add4/Add1/_14_ ));
 OAI21_X2 \Add1/Add4/Add1/_30_  (.A(\Add1/Add4/Add1/_00_ ),
    .B1(\Add1/Add4/Add1/_12_ ),
    .B2(\Add1/Add4/Add1/_13_ ),
    .ZN(\Add1/Add4/c1 ));
 XNOR2_X1 \Add1/Add4/Add1/_31_  (.A(\Add1/c3 ),
    .B(\Add1/Add4/Add1/_05_ ),
    .ZN(s[24]));
 XNOR2_X1 \Add1/Add4/Add1/_32_  (.A(\Add1/Add4/Add1/_06_ ),
    .B(\Add1/Add4/Add1/_08_ ),
    .ZN(s[25]));
 XNOR2_X1 \Add1/Add4/Add1/_33_  (.A(\Add1/Add4/Add1/_09_ ),
    .B(\Add1/Add4/Add1/_11_ ),
    .ZN(s[26]));
 XNOR2_X1 \Add1/Add4/Add1/_34_  (.A(\Add1/Add4/Add1/_12_ ),
    .B(\Add1/Add4/Add1/_14_ ),
    .ZN(s[27]));
 NAND2_X1 \Add1/Add4/Add2/_15_  (.A1(a[31]),
    .A2(b[31]),
    .ZN(\Add1/Add4/Add2/_00_ ));
 AND2_X1 \Add1/Add4/Add2/_16_  (.A1(a[30]),
    .A2(b[30]),
    .ZN(\Add1/Add4/Add2/_01_ ));
 NAND2_X1 \Add1/Add4/Add2/_17_  (.A1(a[29]),
    .A2(b[29]),
    .ZN(\Add1/Add4/Add2/_02_ ));
 AND2_X1 \Add1/Add4/Add2/_18_  (.A1(a[28]),
    .A2(b[28]),
    .ZN(\Add1/Add4/Add2/_03_ ));
 OR2_X1 \Add1/Add4/Add2/_19_  (.A1(a[28]),
    .A2(b[28]),
    .ZN(\Add1/Add4/Add2/_04_ ));
 XNOR2_X1 \Add1/Add4/Add2/_20_  (.A(a[28]),
    .B(b[28]),
    .ZN(\Add1/Add4/Add2/_05_ ));
 AOI21_X2 \Add1/Add4/Add2/_21_  (.A(\Add1/Add4/Add2/_03_ ),
    .B1(\Add1/Add4/Add2/_04_ ),
    .B2(\Add1/Add4/c1 ),
    .ZN(\Add1/Add4/Add2/_06_ ));
 NOR2_X1 \Add1/Add4/Add2/_22_  (.A1(a[29]),
    .A2(b[29]),
    .ZN(\Add1/Add4/Add2/_07_ ));
 XOR2_X1 \Add1/Add4/Add2/_23_  (.A(a[29]),
    .B(b[29]),
    .Z(\Add1/Add4/Add2/_08_ ));
 OAI21_X2 \Add1/Add4/Add2/_24_  (.A(\Add1/Add4/Add2/_02_ ),
    .B1(\Add1/Add4/Add2/_06_ ),
    .B2(\Add1/Add4/Add2/_07_ ),
    .ZN(\Add1/Add4/Add2/_09_ ));
 OR2_X1 \Add1/Add4/Add2/_25_  (.A1(a[30]),
    .A2(b[30]),
    .ZN(\Add1/Add4/Add2/_10_ ));
 XNOR2_X1 \Add1/Add4/Add2/_26_  (.A(a[30]),
    .B(b[30]),
    .ZN(\Add1/Add4/Add2/_11_ ));
 AOI21_X2 \Add1/Add4/Add2/_27_  (.A(\Add1/Add4/Add2/_01_ ),
    .B1(\Add1/Add4/Add2/_09_ ),
    .B2(\Add1/Add4/Add2/_10_ ),
    .ZN(\Add1/Add4/Add2/_12_ ));
 NOR2_X1 \Add1/Add4/Add2/_28_  (.A1(a[31]),
    .A2(b[31]),
    .ZN(\Add1/Add4/Add2/_13_ ));
 XOR2_X1 \Add1/Add4/Add2/_29_  (.A(a[31]),
    .B(b[31]),
    .Z(\Add1/Add4/Add2/_14_ ));
 OAI21_X2 \Add1/Add4/Add2/_30_  (.A(\Add1/Add4/Add2/_00_ ),
    .B1(\Add1/Add4/Add2/_12_ ),
    .B2(\Add1/Add4/Add2/_13_ ),
    .ZN(c1));
 XNOR2_X1 \Add1/Add4/Add2/_31_  (.A(\Add1/Add4/c1 ),
    .B(\Add1/Add4/Add2/_05_ ),
    .ZN(s[28]));
 XNOR2_X1 \Add1/Add4/Add2/_32_  (.A(\Add1/Add4/Add2/_06_ ),
    .B(\Add1/Add4/Add2/_08_ ),
    .ZN(s[29]));
 XNOR2_X1 \Add1/Add4/Add2/_33_  (.A(\Add1/Add4/Add2/_09_ ),
    .B(\Add1/Add4/Add2/_11_ ),
    .ZN(s[30]));
 XNOR2_X1 \Add1/Add4/Add2/_34_  (.A(\Add1/Add4/Add2/_12_ ),
    .B(\Add1/Add4/Add2/_14_ ),
    .ZN(s[31]));
 NAND2_X1 \Add2/Add1/Add1/_15_  (.A1(a[35]),
    .A2(b[35]),
    .ZN(\Add2/Add1/Add1/_00_ ));
 AND2_X1 \Add2/Add1/Add1/_16_  (.A1(a[34]),
    .A2(b[34]),
    .ZN(\Add2/Add1/Add1/_01_ ));
 NAND2_X1 \Add2/Add1/Add1/_17_  (.A1(a[33]),
    .A2(b[33]),
    .ZN(\Add2/Add1/Add1/_02_ ));
 AND2_X1 \Add2/Add1/Add1/_18_  (.A1(a[32]),
    .A2(b[32]),
    .ZN(\Add2/Add1/Add1/_03_ ));
 OR2_X1 \Add2/Add1/Add1/_19_  (.A1(a[32]),
    .A2(b[32]),
    .ZN(\Add2/Add1/Add1/_04_ ));
 XNOR2_X1 \Add2/Add1/Add1/_20_  (.A(a[32]),
    .B(b[32]),
    .ZN(\Add2/Add1/Add1/_05_ ));
 AOI21_X2 \Add2/Add1/Add1/_21_  (.A(\Add2/Add1/Add1/_03_ ),
    .B1(\Add2/Add1/Add1/_04_ ),
    .B2(c1),
    .ZN(\Add2/Add1/Add1/_06_ ));
 NOR2_X1 \Add2/Add1/Add1/_22_  (.A1(a[33]),
    .A2(b[33]),
    .ZN(\Add2/Add1/Add1/_07_ ));
 XOR2_X1 \Add2/Add1/Add1/_23_  (.A(a[33]),
    .B(b[33]),
    .Z(\Add2/Add1/Add1/_08_ ));
 OAI21_X2 \Add2/Add1/Add1/_24_  (.A(\Add2/Add1/Add1/_02_ ),
    .B1(\Add2/Add1/Add1/_06_ ),
    .B2(\Add2/Add1/Add1/_07_ ),
    .ZN(\Add2/Add1/Add1/_09_ ));
 OR2_X1 \Add2/Add1/Add1/_25_  (.A1(a[34]),
    .A2(b[34]),
    .ZN(\Add2/Add1/Add1/_10_ ));
 XNOR2_X1 \Add2/Add1/Add1/_26_  (.A(a[34]),
    .B(b[34]),
    .ZN(\Add2/Add1/Add1/_11_ ));
 AOI21_X2 \Add2/Add1/Add1/_27_  (.A(\Add2/Add1/Add1/_01_ ),
    .B1(\Add2/Add1/Add1/_09_ ),
    .B2(\Add2/Add1/Add1/_10_ ),
    .ZN(\Add2/Add1/Add1/_12_ ));
 NOR2_X1 \Add2/Add1/Add1/_28_  (.A1(a[35]),
    .A2(b[35]),
    .ZN(\Add2/Add1/Add1/_13_ ));
 XOR2_X1 \Add2/Add1/Add1/_29_  (.A(a[35]),
    .B(b[35]),
    .Z(\Add2/Add1/Add1/_14_ ));
 OAI21_X2 \Add2/Add1/Add1/_30_  (.A(\Add2/Add1/Add1/_00_ ),
    .B1(\Add2/Add1/Add1/_12_ ),
    .B2(\Add2/Add1/Add1/_13_ ),
    .ZN(\Add2/Add1/c1 ));
 XNOR2_X1 \Add2/Add1/Add1/_31_  (.A(c1),
    .B(\Add2/Add1/Add1/_05_ ),
    .ZN(s[32]));
 XNOR2_X1 \Add2/Add1/Add1/_32_  (.A(\Add2/Add1/Add1/_06_ ),
    .B(\Add2/Add1/Add1/_08_ ),
    .ZN(s[33]));
 XNOR2_X1 \Add2/Add1/Add1/_33_  (.A(\Add2/Add1/Add1/_09_ ),
    .B(\Add2/Add1/Add1/_11_ ),
    .ZN(s[34]));
 XNOR2_X1 \Add2/Add1/Add1/_34_  (.A(\Add2/Add1/Add1/_12_ ),
    .B(\Add2/Add1/Add1/_14_ ),
    .ZN(s[35]));
 NAND2_X1 \Add2/Add1/Add2/_15_  (.A1(a[39]),
    .A2(b[39]),
    .ZN(\Add2/Add1/Add2/_00_ ));
 AND2_X1 \Add2/Add1/Add2/_16_  (.A1(a[38]),
    .A2(b[38]),
    .ZN(\Add2/Add1/Add2/_01_ ));
 NAND2_X1 \Add2/Add1/Add2/_17_  (.A1(a[37]),
    .A2(b[37]),
    .ZN(\Add2/Add1/Add2/_02_ ));
 AND2_X1 \Add2/Add1/Add2/_18_  (.A1(a[36]),
    .A2(b[36]),
    .ZN(\Add2/Add1/Add2/_03_ ));
 OR2_X1 \Add2/Add1/Add2/_19_  (.A1(a[36]),
    .A2(b[36]),
    .ZN(\Add2/Add1/Add2/_04_ ));
 XNOR2_X1 \Add2/Add1/Add2/_20_  (.A(a[36]),
    .B(b[36]),
    .ZN(\Add2/Add1/Add2/_05_ ));
 AOI21_X2 \Add2/Add1/Add2/_21_  (.A(\Add2/Add1/Add2/_03_ ),
    .B1(\Add2/Add1/Add2/_04_ ),
    .B2(\Add2/Add1/c1 ),
    .ZN(\Add2/Add1/Add2/_06_ ));
 NOR2_X1 \Add2/Add1/Add2/_22_  (.A1(a[37]),
    .A2(b[37]),
    .ZN(\Add2/Add1/Add2/_07_ ));
 XOR2_X1 \Add2/Add1/Add2/_23_  (.A(a[37]),
    .B(b[37]),
    .Z(\Add2/Add1/Add2/_08_ ));
 OAI21_X2 \Add2/Add1/Add2/_24_  (.A(\Add2/Add1/Add2/_02_ ),
    .B1(\Add2/Add1/Add2/_06_ ),
    .B2(\Add2/Add1/Add2/_07_ ),
    .ZN(\Add2/Add1/Add2/_09_ ));
 OR2_X1 \Add2/Add1/Add2/_25_  (.A1(a[38]),
    .A2(b[38]),
    .ZN(\Add2/Add1/Add2/_10_ ));
 XNOR2_X1 \Add2/Add1/Add2/_26_  (.A(a[38]),
    .B(b[38]),
    .ZN(\Add2/Add1/Add2/_11_ ));
 AOI21_X2 \Add2/Add1/Add2/_27_  (.A(\Add2/Add1/Add2/_01_ ),
    .B1(\Add2/Add1/Add2/_09_ ),
    .B2(\Add2/Add1/Add2/_10_ ),
    .ZN(\Add2/Add1/Add2/_12_ ));
 NOR2_X1 \Add2/Add1/Add2/_28_  (.A1(a[39]),
    .A2(b[39]),
    .ZN(\Add2/Add1/Add2/_13_ ));
 XOR2_X1 \Add2/Add1/Add2/_29_  (.A(a[39]),
    .B(b[39]),
    .Z(\Add2/Add1/Add2/_14_ ));
 OAI21_X2 \Add2/Add1/Add2/_30_  (.A(\Add2/Add1/Add2/_00_ ),
    .B1(\Add2/Add1/Add2/_12_ ),
    .B2(\Add2/Add1/Add2/_13_ ),
    .ZN(\Add2/c1 ));
 XNOR2_X1 \Add2/Add1/Add2/_31_  (.A(\Add2/Add1/c1 ),
    .B(\Add2/Add1/Add2/_05_ ),
    .ZN(s[36]));
 XNOR2_X1 \Add2/Add1/Add2/_32_  (.A(\Add2/Add1/Add2/_06_ ),
    .B(\Add2/Add1/Add2/_08_ ),
    .ZN(s[37]));
 XNOR2_X1 \Add2/Add1/Add2/_33_  (.A(\Add2/Add1/Add2/_09_ ),
    .B(\Add2/Add1/Add2/_11_ ),
    .ZN(s[38]));
 XNOR2_X1 \Add2/Add1/Add2/_34_  (.A(\Add2/Add1/Add2/_12_ ),
    .B(\Add2/Add1/Add2/_14_ ),
    .ZN(s[39]));
 NAND2_X1 \Add2/Add2/Add1/_15_  (.A1(a[43]),
    .A2(b[43]),
    .ZN(\Add2/Add2/Add1/_00_ ));
 AND2_X1 \Add2/Add2/Add1/_16_  (.A1(a[42]),
    .A2(b[42]),
    .ZN(\Add2/Add2/Add1/_01_ ));
 NAND2_X1 \Add2/Add2/Add1/_17_  (.A1(a[41]),
    .A2(b[41]),
    .ZN(\Add2/Add2/Add1/_02_ ));
 AND2_X1 \Add2/Add2/Add1/_18_  (.A1(a[40]),
    .A2(b[40]),
    .ZN(\Add2/Add2/Add1/_03_ ));
 OR2_X1 \Add2/Add2/Add1/_19_  (.A1(a[40]),
    .A2(b[40]),
    .ZN(\Add2/Add2/Add1/_04_ ));
 XNOR2_X1 \Add2/Add2/Add1/_20_  (.A(a[40]),
    .B(b[40]),
    .ZN(\Add2/Add2/Add1/_05_ ));
 AOI21_X2 \Add2/Add2/Add1/_21_  (.A(\Add2/Add2/Add1/_03_ ),
    .B1(\Add2/Add2/Add1/_04_ ),
    .B2(\Add2/c1 ),
    .ZN(\Add2/Add2/Add1/_06_ ));
 NOR2_X1 \Add2/Add2/Add1/_22_  (.A1(a[41]),
    .A2(b[41]),
    .ZN(\Add2/Add2/Add1/_07_ ));
 XOR2_X1 \Add2/Add2/Add1/_23_  (.A(a[41]),
    .B(b[41]),
    .Z(\Add2/Add2/Add1/_08_ ));
 OAI21_X1 \Add2/Add2/Add1/_24_  (.A(\Add2/Add2/Add1/_02_ ),
    .B1(\Add2/Add2/Add1/_06_ ),
    .B2(\Add2/Add2/Add1/_07_ ),
    .ZN(\Add2/Add2/Add1/_09_ ));
 OR2_X1 \Add2/Add2/Add1/_25_  (.A1(a[42]),
    .A2(b[42]),
    .ZN(\Add2/Add2/Add1/_10_ ));
 XNOR2_X1 \Add2/Add2/Add1/_26_  (.A(a[42]),
    .B(b[42]),
    .ZN(\Add2/Add2/Add1/_11_ ));
 AOI21_X2 \Add2/Add2/Add1/_27_  (.A(\Add2/Add2/Add1/_01_ ),
    .B1(\Add2/Add2/Add1/_09_ ),
    .B2(\Add2/Add2/Add1/_10_ ),
    .ZN(\Add2/Add2/Add1/_12_ ));
 NOR2_X1 \Add2/Add2/Add1/_28_  (.A1(a[43]),
    .A2(b[43]),
    .ZN(\Add2/Add2/Add1/_13_ ));
 XOR2_X1 \Add2/Add2/Add1/_29_  (.A(a[43]),
    .B(b[43]),
    .Z(\Add2/Add2/Add1/_14_ ));
 OAI21_X2 \Add2/Add2/Add1/_30_  (.A(\Add2/Add2/Add1/_00_ ),
    .B1(\Add2/Add2/Add1/_12_ ),
    .B2(\Add2/Add2/Add1/_13_ ),
    .ZN(\Add2/Add2/c1 ));
 XNOR2_X1 \Add2/Add2/Add1/_31_  (.A(\Add2/c1 ),
    .B(\Add2/Add2/Add1/_05_ ),
    .ZN(s[40]));
 XNOR2_X1 \Add2/Add2/Add1/_32_  (.A(\Add2/Add2/Add1/_06_ ),
    .B(\Add2/Add2/Add1/_08_ ),
    .ZN(s[41]));
 XNOR2_X1 \Add2/Add2/Add1/_33_  (.A(\Add2/Add2/Add1/_09_ ),
    .B(\Add2/Add2/Add1/_11_ ),
    .ZN(s[42]));
 XNOR2_X1 \Add2/Add2/Add1/_34_  (.A(\Add2/Add2/Add1/_12_ ),
    .B(\Add2/Add2/Add1/_14_ ),
    .ZN(s[43]));
 NAND2_X1 \Add2/Add2/Add2/_15_  (.A1(a[47]),
    .A2(b[47]),
    .ZN(\Add2/Add2/Add2/_00_ ));
 AND2_X1 \Add2/Add2/Add2/_16_  (.A1(a[46]),
    .A2(b[46]),
    .ZN(\Add2/Add2/Add2/_01_ ));
 NAND2_X1 \Add2/Add2/Add2/_17_  (.A1(a[45]),
    .A2(b[45]),
    .ZN(\Add2/Add2/Add2/_02_ ));
 AND2_X1 \Add2/Add2/Add2/_18_  (.A1(a[44]),
    .A2(b[44]),
    .ZN(\Add2/Add2/Add2/_03_ ));
 OR2_X1 \Add2/Add2/Add2/_19_  (.A1(a[44]),
    .A2(b[44]),
    .ZN(\Add2/Add2/Add2/_04_ ));
 XNOR2_X1 \Add2/Add2/Add2/_20_  (.A(a[44]),
    .B(b[44]),
    .ZN(\Add2/Add2/Add2/_05_ ));
 AOI21_X2 \Add2/Add2/Add2/_21_  (.A(\Add2/Add2/Add2/_03_ ),
    .B1(\Add2/Add2/Add2/_04_ ),
    .B2(\Add2/Add2/c1 ),
    .ZN(\Add2/Add2/Add2/_06_ ));
 NOR2_X1 \Add2/Add2/Add2/_22_  (.A1(a[45]),
    .A2(b[45]),
    .ZN(\Add2/Add2/Add2/_07_ ));
 XOR2_X1 \Add2/Add2/Add2/_23_  (.A(a[45]),
    .B(b[45]),
    .Z(\Add2/Add2/Add2/_08_ ));
 OAI21_X2 \Add2/Add2/Add2/_24_  (.A(\Add2/Add2/Add2/_02_ ),
    .B1(\Add2/Add2/Add2/_06_ ),
    .B2(\Add2/Add2/Add2/_07_ ),
    .ZN(\Add2/Add2/Add2/_09_ ));
 OR2_X1 \Add2/Add2/Add2/_25_  (.A1(a[46]),
    .A2(b[46]),
    .ZN(\Add2/Add2/Add2/_10_ ));
 XNOR2_X1 \Add2/Add2/Add2/_26_  (.A(a[46]),
    .B(b[46]),
    .ZN(\Add2/Add2/Add2/_11_ ));
 AOI21_X2 \Add2/Add2/Add2/_27_  (.A(\Add2/Add2/Add2/_01_ ),
    .B1(\Add2/Add2/Add2/_09_ ),
    .B2(\Add2/Add2/Add2/_10_ ),
    .ZN(\Add2/Add2/Add2/_12_ ));
 NOR2_X1 \Add2/Add2/Add2/_28_  (.A1(a[47]),
    .A2(b[47]),
    .ZN(\Add2/Add2/Add2/_13_ ));
 XOR2_X1 \Add2/Add2/Add2/_29_  (.A(a[47]),
    .B(b[47]),
    .Z(\Add2/Add2/Add2/_14_ ));
 OAI21_X2 \Add2/Add2/Add2/_30_  (.A(\Add2/Add2/Add2/_00_ ),
    .B1(\Add2/Add2/Add2/_12_ ),
    .B2(\Add2/Add2/Add2/_13_ ),
    .ZN(\Add2/c2 ));
 XNOR2_X1 \Add2/Add2/Add2/_31_  (.A(\Add2/Add2/c1 ),
    .B(\Add2/Add2/Add2/_05_ ),
    .ZN(s[44]));
 XNOR2_X1 \Add2/Add2/Add2/_32_  (.A(\Add2/Add2/Add2/_06_ ),
    .B(\Add2/Add2/Add2/_08_ ),
    .ZN(s[45]));
 XNOR2_X1 \Add2/Add2/Add2/_33_  (.A(\Add2/Add2/Add2/_09_ ),
    .B(\Add2/Add2/Add2/_11_ ),
    .ZN(s[46]));
 XNOR2_X1 \Add2/Add2/Add2/_34_  (.A(\Add2/Add2/Add2/_12_ ),
    .B(\Add2/Add2/Add2/_14_ ),
    .ZN(s[47]));
 NAND2_X1 \Add2/Add3/Add1/_15_  (.A1(a[51]),
    .A2(b[51]),
    .ZN(\Add2/Add3/Add1/_00_ ));
 AND2_X1 \Add2/Add3/Add1/_16_  (.A1(a[50]),
    .A2(b[50]),
    .ZN(\Add2/Add3/Add1/_01_ ));
 NAND2_X1 \Add2/Add3/Add1/_17_  (.A1(a[49]),
    .A2(b[49]),
    .ZN(\Add2/Add3/Add1/_02_ ));
 AND2_X1 \Add2/Add3/Add1/_18_  (.A1(a[48]),
    .A2(b[48]),
    .ZN(\Add2/Add3/Add1/_03_ ));
 OR2_X1 \Add2/Add3/Add1/_19_  (.A1(a[48]),
    .A2(b[48]),
    .ZN(\Add2/Add3/Add1/_04_ ));
 XNOR2_X1 \Add2/Add3/Add1/_20_  (.A(a[48]),
    .B(b[48]),
    .ZN(\Add2/Add3/Add1/_05_ ));
 AOI21_X2 \Add2/Add3/Add1/_21_  (.A(\Add2/Add3/Add1/_03_ ),
    .B1(\Add2/Add3/Add1/_04_ ),
    .B2(\Add2/c2 ),
    .ZN(\Add2/Add3/Add1/_06_ ));
 NOR2_X1 \Add2/Add3/Add1/_22_  (.A1(a[49]),
    .A2(b[49]),
    .ZN(\Add2/Add3/Add1/_07_ ));
 XOR2_X1 \Add2/Add3/Add1/_23_  (.A(a[49]),
    .B(b[49]),
    .Z(\Add2/Add3/Add1/_08_ ));
 OAI21_X2 \Add2/Add3/Add1/_24_  (.A(\Add2/Add3/Add1/_02_ ),
    .B1(\Add2/Add3/Add1/_06_ ),
    .B2(\Add2/Add3/Add1/_07_ ),
    .ZN(\Add2/Add3/Add1/_09_ ));
 OR2_X1 \Add2/Add3/Add1/_25_  (.A1(a[50]),
    .A2(b[50]),
    .ZN(\Add2/Add3/Add1/_10_ ));
 XNOR2_X1 \Add2/Add3/Add1/_26_  (.A(a[50]),
    .B(b[50]),
    .ZN(\Add2/Add3/Add1/_11_ ));
 AOI21_X2 \Add2/Add3/Add1/_27_  (.A(\Add2/Add3/Add1/_01_ ),
    .B1(\Add2/Add3/Add1/_09_ ),
    .B2(\Add2/Add3/Add1/_10_ ),
    .ZN(\Add2/Add3/Add1/_12_ ));
 NOR2_X1 \Add2/Add3/Add1/_28_  (.A1(a[51]),
    .A2(b[51]),
    .ZN(\Add2/Add3/Add1/_13_ ));
 XOR2_X1 \Add2/Add3/Add1/_29_  (.A(a[51]),
    .B(b[51]),
    .Z(\Add2/Add3/Add1/_14_ ));
 OAI21_X2 \Add2/Add3/Add1/_30_  (.A(\Add2/Add3/Add1/_00_ ),
    .B1(\Add2/Add3/Add1/_12_ ),
    .B2(\Add2/Add3/Add1/_13_ ),
    .ZN(\Add2/Add3/c1 ));
 XNOR2_X1 \Add2/Add3/Add1/_31_  (.A(\Add2/c2 ),
    .B(\Add2/Add3/Add1/_05_ ),
    .ZN(s[48]));
 XNOR2_X1 \Add2/Add3/Add1/_32_  (.A(\Add2/Add3/Add1/_06_ ),
    .B(\Add2/Add3/Add1/_08_ ),
    .ZN(s[49]));
 XNOR2_X1 \Add2/Add3/Add1/_33_  (.A(\Add2/Add3/Add1/_09_ ),
    .B(\Add2/Add3/Add1/_11_ ),
    .ZN(s[50]));
 XNOR2_X1 \Add2/Add3/Add1/_34_  (.A(\Add2/Add3/Add1/_12_ ),
    .B(\Add2/Add3/Add1/_14_ ),
    .ZN(s[51]));
 NAND2_X1 \Add2/Add3/Add2/_15_  (.A1(a[55]),
    .A2(b[55]),
    .ZN(\Add2/Add3/Add2/_00_ ));
 AND2_X1 \Add2/Add3/Add2/_16_  (.A1(a[54]),
    .A2(b[54]),
    .ZN(\Add2/Add3/Add2/_01_ ));
 NAND2_X1 \Add2/Add3/Add2/_17_  (.A1(a[53]),
    .A2(b[53]),
    .ZN(\Add2/Add3/Add2/_02_ ));
 AND2_X1 \Add2/Add3/Add2/_18_  (.A1(a[52]),
    .A2(b[52]),
    .ZN(\Add2/Add3/Add2/_03_ ));
 OR2_X1 \Add2/Add3/Add2/_19_  (.A1(a[52]),
    .A2(b[52]),
    .ZN(\Add2/Add3/Add2/_04_ ));
 XNOR2_X1 \Add2/Add3/Add2/_20_  (.A(a[52]),
    .B(b[52]),
    .ZN(\Add2/Add3/Add2/_05_ ));
 AOI21_X2 \Add2/Add3/Add2/_21_  (.A(\Add2/Add3/Add2/_03_ ),
    .B1(\Add2/Add3/Add2/_04_ ),
    .B2(\Add2/Add3/c1 ),
    .ZN(\Add2/Add3/Add2/_06_ ));
 NOR2_X1 \Add2/Add3/Add2/_22_  (.A1(a[53]),
    .A2(b[53]),
    .ZN(\Add2/Add3/Add2/_07_ ));
 XOR2_X1 \Add2/Add3/Add2/_23_  (.A(a[53]),
    .B(b[53]),
    .Z(\Add2/Add3/Add2/_08_ ));
 OAI21_X1 \Add2/Add3/Add2/_24_  (.A(\Add2/Add3/Add2/_02_ ),
    .B1(\Add2/Add3/Add2/_06_ ),
    .B2(\Add2/Add3/Add2/_07_ ),
    .ZN(\Add2/Add3/Add2/_09_ ));
 OR2_X1 \Add2/Add3/Add2/_25_  (.A1(a[54]),
    .A2(b[54]),
    .ZN(\Add2/Add3/Add2/_10_ ));
 XNOR2_X1 \Add2/Add3/Add2/_26_  (.A(a[54]),
    .B(b[54]),
    .ZN(\Add2/Add3/Add2/_11_ ));
 AOI21_X2 \Add2/Add3/Add2/_27_  (.A(\Add2/Add3/Add2/_01_ ),
    .B1(\Add2/Add3/Add2/_09_ ),
    .B2(\Add2/Add3/Add2/_10_ ),
    .ZN(\Add2/Add3/Add2/_12_ ));
 NOR2_X1 \Add2/Add3/Add2/_28_  (.A1(a[55]),
    .A2(b[55]),
    .ZN(\Add2/Add3/Add2/_13_ ));
 XOR2_X1 \Add2/Add3/Add2/_29_  (.A(a[55]),
    .B(b[55]),
    .Z(\Add2/Add3/Add2/_14_ ));
 OAI21_X2 \Add2/Add3/Add2/_30_  (.A(\Add2/Add3/Add2/_00_ ),
    .B1(\Add2/Add3/Add2/_12_ ),
    .B2(\Add2/Add3/Add2/_13_ ),
    .ZN(\Add2/c3 ));
 XNOR2_X1 \Add2/Add3/Add2/_31_  (.A(\Add2/Add3/c1 ),
    .B(\Add2/Add3/Add2/_05_ ),
    .ZN(s[52]));
 XNOR2_X1 \Add2/Add3/Add2/_32_  (.A(\Add2/Add3/Add2/_06_ ),
    .B(\Add2/Add3/Add2/_08_ ),
    .ZN(s[53]));
 XNOR2_X1 \Add2/Add3/Add2/_33_  (.A(\Add2/Add3/Add2/_09_ ),
    .B(\Add2/Add3/Add2/_11_ ),
    .ZN(s[54]));
 XNOR2_X1 \Add2/Add3/Add2/_34_  (.A(\Add2/Add3/Add2/_12_ ),
    .B(\Add2/Add3/Add2/_14_ ),
    .ZN(s[55]));
 NAND2_X1 \Add2/Add4/Add1/_15_  (.A1(a[59]),
    .A2(b[59]),
    .ZN(\Add2/Add4/Add1/_00_ ));
 AND2_X1 \Add2/Add4/Add1/_16_  (.A1(a[58]),
    .A2(b[58]),
    .ZN(\Add2/Add4/Add1/_01_ ));
 NAND2_X1 \Add2/Add4/Add1/_17_  (.A1(a[57]),
    .A2(b[57]),
    .ZN(\Add2/Add4/Add1/_02_ ));
 AND2_X1 \Add2/Add4/Add1/_18_  (.A1(a[56]),
    .A2(b[56]),
    .ZN(\Add2/Add4/Add1/_03_ ));
 OR2_X1 \Add2/Add4/Add1/_19_  (.A1(a[56]),
    .A2(b[56]),
    .ZN(\Add2/Add4/Add1/_04_ ));
 XNOR2_X1 \Add2/Add4/Add1/_20_  (.A(a[56]),
    .B(b[56]),
    .ZN(\Add2/Add4/Add1/_05_ ));
 AOI21_X2 \Add2/Add4/Add1/_21_  (.A(\Add2/Add4/Add1/_03_ ),
    .B1(\Add2/Add4/Add1/_04_ ),
    .B2(\Add2/c3 ),
    .ZN(\Add2/Add4/Add1/_06_ ));
 NOR2_X1 \Add2/Add4/Add1/_22_  (.A1(a[57]),
    .A2(b[57]),
    .ZN(\Add2/Add4/Add1/_07_ ));
 XOR2_X1 \Add2/Add4/Add1/_23_  (.A(a[57]),
    .B(b[57]),
    .Z(\Add2/Add4/Add1/_08_ ));
 OAI21_X2 \Add2/Add4/Add1/_24_  (.A(\Add2/Add4/Add1/_02_ ),
    .B1(\Add2/Add4/Add1/_06_ ),
    .B2(\Add2/Add4/Add1/_07_ ),
    .ZN(\Add2/Add4/Add1/_09_ ));
 OR2_X1 \Add2/Add4/Add1/_25_  (.A1(a[58]),
    .A2(b[58]),
    .ZN(\Add2/Add4/Add1/_10_ ));
 XNOR2_X1 \Add2/Add4/Add1/_26_  (.A(a[58]),
    .B(b[58]),
    .ZN(\Add2/Add4/Add1/_11_ ));
 AOI21_X2 \Add2/Add4/Add1/_27_  (.A(\Add2/Add4/Add1/_01_ ),
    .B1(\Add2/Add4/Add1/_09_ ),
    .B2(\Add2/Add4/Add1/_10_ ),
    .ZN(\Add2/Add4/Add1/_12_ ));
 NOR2_X1 \Add2/Add4/Add1/_28_  (.A1(a[59]),
    .A2(b[59]),
    .ZN(\Add2/Add4/Add1/_13_ ));
 XOR2_X1 \Add2/Add4/Add1/_29_  (.A(a[59]),
    .B(b[59]),
    .Z(\Add2/Add4/Add1/_14_ ));
 OAI21_X2 \Add2/Add4/Add1/_30_  (.A(\Add2/Add4/Add1/_00_ ),
    .B1(\Add2/Add4/Add1/_12_ ),
    .B2(\Add2/Add4/Add1/_13_ ),
    .ZN(\Add2/Add4/c1 ));
 XNOR2_X1 \Add2/Add4/Add1/_31_  (.A(\Add2/c3 ),
    .B(\Add2/Add4/Add1/_05_ ),
    .ZN(s[56]));
 XNOR2_X1 \Add2/Add4/Add1/_32_  (.A(\Add2/Add4/Add1/_06_ ),
    .B(\Add2/Add4/Add1/_08_ ),
    .ZN(s[57]));
 XNOR2_X1 \Add2/Add4/Add1/_33_  (.A(\Add2/Add4/Add1/_09_ ),
    .B(\Add2/Add4/Add1/_11_ ),
    .ZN(s[58]));
 XNOR2_X1 \Add2/Add4/Add1/_34_  (.A(\Add2/Add4/Add1/_12_ ),
    .B(\Add2/Add4/Add1/_14_ ),
    .ZN(s[59]));
 NAND2_X1 \Add2/Add4/Add2/_15_  (.A1(a[63]),
    .A2(b[63]),
    .ZN(\Add2/Add4/Add2/_00_ ));
 AND2_X1 \Add2/Add4/Add2/_16_  (.A1(a[62]),
    .A2(b[62]),
    .ZN(\Add2/Add4/Add2/_01_ ));
 NAND2_X1 \Add2/Add4/Add2/_17_  (.A1(a[61]),
    .A2(b[61]),
    .ZN(\Add2/Add4/Add2/_02_ ));
 AND2_X1 \Add2/Add4/Add2/_18_  (.A1(a[60]),
    .A2(b[60]),
    .ZN(\Add2/Add4/Add2/_03_ ));
 OR2_X1 \Add2/Add4/Add2/_19_  (.A1(a[60]),
    .A2(b[60]),
    .ZN(\Add2/Add4/Add2/_04_ ));
 XNOR2_X1 \Add2/Add4/Add2/_20_  (.A(a[60]),
    .B(b[60]),
    .ZN(\Add2/Add4/Add2/_05_ ));
 AOI21_X2 \Add2/Add4/Add2/_21_  (.A(\Add2/Add4/Add2/_03_ ),
    .B1(\Add2/Add4/Add2/_04_ ),
    .B2(\Add2/Add4/c1 ),
    .ZN(\Add2/Add4/Add2/_06_ ));
 NOR2_X1 \Add2/Add4/Add2/_22_  (.A1(a[61]),
    .A2(b[61]),
    .ZN(\Add2/Add4/Add2/_07_ ));
 XOR2_X1 \Add2/Add4/Add2/_23_  (.A(a[61]),
    .B(b[61]),
    .Z(\Add2/Add4/Add2/_08_ ));
 OAI21_X2 \Add2/Add4/Add2/_24_  (.A(\Add2/Add4/Add2/_02_ ),
    .B1(\Add2/Add4/Add2/_06_ ),
    .B2(\Add2/Add4/Add2/_07_ ),
    .ZN(\Add2/Add4/Add2/_09_ ));
 OR2_X1 \Add2/Add4/Add2/_25_  (.A1(a[62]),
    .A2(b[62]),
    .ZN(\Add2/Add4/Add2/_10_ ));
 XNOR2_X1 \Add2/Add4/Add2/_26_  (.A(a[62]),
    .B(b[62]),
    .ZN(\Add2/Add4/Add2/_11_ ));
 AOI21_X1 \Add2/Add4/Add2/_27_  (.A(\Add2/Add4/Add2/_01_ ),
    .B1(\Add2/Add4/Add2/_09_ ),
    .B2(\Add2/Add4/Add2/_10_ ),
    .ZN(\Add2/Add4/Add2/_12_ ));
 NOR2_X1 \Add2/Add4/Add2/_28_  (.A1(a[63]),
    .A2(b[63]),
    .ZN(\Add2/Add4/Add2/_13_ ));
 XOR2_X1 \Add2/Add4/Add2/_29_  (.A(a[63]),
    .B(b[63]),
    .Z(\Add2/Add4/Add2/_14_ ));
 OAI21_X1 \Add2/Add4/Add2/_30_  (.A(\Add2/Add4/Add2/_00_ ),
    .B1(\Add2/Add4/Add2/_12_ ),
    .B2(\Add2/Add4/Add2/_13_ ),
    .ZN(cout));
 XNOR2_X1 \Add2/Add4/Add2/_31_  (.A(\Add2/Add4/c1 ),
    .B(\Add2/Add4/Add2/_05_ ),
    .ZN(s[60]));
 XNOR2_X1 \Add2/Add4/Add2/_32_  (.A(\Add2/Add4/Add2/_06_ ),
    .B(\Add2/Add4/Add2/_08_ ),
    .ZN(s[61]));
 XNOR2_X1 \Add2/Add4/Add2/_33_  (.A(\Add2/Add4/Add2/_09_ ),
    .B(\Add2/Add4/Add2/_11_ ),
    .ZN(s[62]));
 XNOR2_X1 \Add2/Add4/Add2/_34_  (.A(\Add2/Add4/Add2/_12_ ),
    .B(\Add2/Add4/Add2/_14_ ),
    .ZN(s[63]));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_113 ();
endmodule
